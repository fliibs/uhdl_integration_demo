module axi_slave #(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 32,
	parameter ID_WIDTH   = 7,
	parameter USER_WIDTH = 5

)(		
		input                   clk,
        input                   rst_n,
		input    [ADDR_WIDTH-1 : 0]                  s0_axi_awaddr,
		input    [2 : 0]                             s0_axi_awprot,
		input                                        s0_axi_awvalid,
		output                                       s0_axi_awready,
		input    [DATA_WIDTH-1 : 0]                  s0_axi_wdata,
		input    [DATA_WIDTH/8-1 : 0]              	 s0_axi_wstrb,
		input                                        s0_axi_wvalid,
		output                                       s0_axi_wready,
		output   [1 : 0]                             s0_axi_bresp,
		output                                       s0_axi_bvalid,
		input                                        s0_axi_bready,
		input    [ADDR_WIDTH-1 : 0]                  s0_axi_araddr,
		input    [2 : 0]                             s0_axi_arprot,
		input                                        s0_axi_arvalid,
		output                                       s0_axi_arready,
		output   [DATA_WIDTH-1 : 0]                  s0_axi_rdata,
		output   [1 : 0]                             s0_axi_rresp,
		output                                       s0_axi_rvalid,
		input                                        s0_axi_rready,

		input   [ID_WIDTH-1 : 0]                       s_axi_awid,
		input   [ADDR_WIDTH-1 : 0]                     s_axi_awaddr,
		input   [7 : 0]                                s_axi_awlen,
		input   [2 : 0]                                s_axi_awsize,
		input   [1 : 0]                                s_axi_awburst,
		input                                          s_axi_awlock,
		input   [3 : 0]                                s_axi_awcache,
		input   [2 : 0]                                s_axi_awprot,
		input   [3 : 0]                                s_axi_awqos,
		input   [USER_WIDTH-1 : 0]                     s_axi_awuser,
		input                                          s_axi_awvalid,
		output                                           s_axi_awready,
		input   [DATA_WIDTH-1 : 0]                     s_axi_wdata,
		input   [DATA_WIDTH/8-1 : 0]                   s_axi_wstrb,
		input                                          s_axi_wlast,
		input   [USER_WIDTH-1 : 0]                     s_axi_wuser,
		input                                          s_axi_wvalid,
		output                                           s_axi_wready,
		output    [ID_WIDTH-1 : 0]                       s_axi_bid,
		output    [1 : 0]                                s_axi_bresp,
		output    [USER_WIDTH-1 : 0]                     s_axi_buser,
		output                                           s_axi_bvalid,
		input                                          s_axi_bready,
		input   [ID_WIDTH-1 : 0]                       s_axi_arid,
		input   [ADDR_WIDTH-1 : 0]                     s_axi_araddr,
		input   [7 : 0]                                s_axi_arlen,
		input   [2 : 0]                                s_axi_arsize,
		input   [1 : 0]                                s_axi_arburst,
		input                                          s_axi_arlock,
		input   [3 : 0]                                s_axi_arcache,
		input   [2 : 0]                                s_axi_arprot,
		input   [3 : 0]                                s_axi_arqos,
		input   [USER_WIDTH-1 : 0]                     s_axi_aruser,
		input    										s_axi_arvalid,
		output     										s_axi_arready,
		output    [ID_WIDTH-1 : 0] 						s_axi_rid,
		output    [DATA_WIDTH-1 : 0] 					s_axi_rdata,
		output    [1 : 0] 								s_axi_rresp,
		output     										s_axi_rlast,
		output    [USER_WIDTH-1 : 0] 					s_axi_ruser,
		output     										s_axi_rvalid,
		input    										s_axi_rready
);


endmodule