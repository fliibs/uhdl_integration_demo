module axi_master #(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 32,
	parameter ID_WIDTH   = 7,
	parameter USER_WIDTH = 5
)(
        input                   clk,
        input                   rst_n,

		output   [ID_WIDTH-1 : 0]                       m_axi_awid,
		output   [ADDR_WIDTH-1 : 0]                     m_axi_awaddr,
		output   [7 : 0]                                m_axi_awlen,
		output   [2 : 0]                                m_axi_awsize,
		output   [1 : 0]                                m_axi_awburst,
		output                                          m_axi_awlock,
		output   [3 : 0]                                m_axi_awcache,
		output   [2 : 0]                                m_axi_awprot,
		output   [3 : 0]                                m_axi_awqos,
		output   [USER_WIDTH-1 : 0]                     m_axi_awuser,
		output                                          m_axi_awvalid,
		input                                           m_axi_awready,
		output   [DATA_WIDTH-1 : 0]                     m_axi_wdata,
		output   [DATA_WIDTH/8-1 : 0]                   m_axi_wstrb,
		output                                          m_axi_wlast,
		output   [USER_WIDTH-1 : 0]                     m_axi_wuser,
		output                                          m_axi_wvalid,
		input                                           m_axi_wready,
		input    [ID_WIDTH-1 : 0]                       m_axi_bid,
		input    [1 : 0]                                m_axi_bresp,
		input    [USER_WIDTH-1 : 0]                     m_axi_buser,
		input                                           m_axi_bvalid,
		output                                          m_axi_bready,
		output   [ID_WIDTH-1 : 0]                       m_axi_arid,
		output   [ADDR_WIDTH-1 : 0]                     m_axi_araddr,
		output   [7 : 0]                                m_axi_arlen,
		output   [2 : 0]                                m_axi_arsize,
		output   [1 : 0]                                m_axi_arburst,
		output                                          m_axi_arlock,
		output   [3 : 0]                                m_axi_arcache,
		output   [2 : 0]                                m_axi_arprot,
		output   [3 : 0]                                m_axi_arqos,
		output   [USER_WIDTH-1 : 0]                     m_axi_aruser,
		output    										m_axi_arvalid,
		input     										m_axi_arready,
		input    [ID_WIDTH-1 : 0] 						m_axi_rid,
		input    [DATA_WIDTH-1 : 0] 					m_axi_rdata,
		input    [1 : 0] 								m_axi_rresp,
		input     										m_axi_rlast,
		input    [USER_WIDTH-1 : 0] 					m_axi_ruser,
		input     										m_axi_rvalid,
		output    										m_axi_rready

);


endmodule