module demo_inout (
    input  data_tri,
    input  data_tx,
    output data_rx,
    inout  data_io_2
  );

endmodule
